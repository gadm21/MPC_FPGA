module model();

endmodule